


`timescale 1ps/1ps
module tb_mul_f();
			parameter msb = 31, T = 2;
			
			reg[msb:0] A, B;
			reg[7:0] S;
			wire[msb:0] O;
			
initial begin
		S = 0;
// === S0 ============
   A = 32'b0_1111111_10000000000000000000000 ;    // 1.5
   B = 32'b0_10000000_00001000000000000000000 ;    // 2.0625
// === S1 ============
#T A = 32'b0_10000000_10000000000000000000000 ;    // 3.0
   B = 32'b0_10000000_11001000000000000000000 ;    // 3.5625
// === S2 ============
#T A = 32'b0_10000001_00100000000000000000000 ;    // 4.5
   B = 32'b0_10000001_01000100000000000000000 ;    // 5.0625
// === S3 ============
#T A = 32'b0_10000001_10000000000000000000000 ;    // 6.0
   B = 32'b0_10000001_10100100000000000000000 ;    // 6.5625
// === S4 ============
#T A = 32'b0_10000001_11100000000000000000000 ;    // 7.5
   B = 32'b0_10000010_00000010000000000000000 ;    // 8.0625
// === S5 ============
#T A = 32'b0_10000010_00100000000000000000000 ;    // 9.0
   B = 32'b0_10000010_00110010000000000000000 ;    // 9.5625
// === S6 ============
#T A = 32'b0_10000010_01010000000000000000000 ;    // 10.5
   B = 32'b0_10000010_01100010000000000000000 ;    // 11.0625
// === S7 ============
#T A = 32'b0_10000010_10000000000000000000000 ;    // 12.0
   B = 32'b0_10000010_10010010000000000000000 ;    // 12.5625
// === S8 ============
#T A = 32'b0_10000010_10110000000000000000000 ;    // 13.5
   B = 32'b0_10000010_11000010000000000000000 ;    // 14.0625
// === S9 ============
#T A = 32'b0_10000010_11100000000000000000000 ;    // 15.0
   B = 32'b0_10000010_11110010000000000000000 ;    // 15.5625
end
			always #T S = S + 1;
			mul_f m(.A(A), .B(B), .O(O));
			
endmodule

